module module_name (input [size] input_name,
                    output [size] output_name);

endmodule