`timescale 1ns / 1ps
//ALU??
module ALU(OP,A,B,F,ZF,CF,OF,SF,PF);
    parameter SIZE = 32;//????
    input [3:0] OP;//????
    input [SIZE:1] A;//????
    input [SIZE:1] B;//????
    output [SIZE:1] F;//????
    output  ZF, //0???, ?????0(??)??1, ???0 
            CF, //??????, ??????C,???C=1?CF=1?????,???C=0?CF=1?????
            OF, //????????????????????OF=1????0
            SF, //???????F??????
            PF; //??????F????1??PF=1????0
    reg [SIZE:1] F;
    reg C,ZF,CF,OF,SF,PF;//C??????
    always@(*)
    begin
        C=0;
        case(OP)
            4'b0000:begin F=A&B; end    //???
            4'b0001:begin F=A|B; end    //???
            4'b0010:begin F=A^B; end    //????
            4'b0011:begin F=~(A|B); end //????
            4'b0100:begin {C,F}=A+B; end //??
            4'b0101:begin {C,F}=A-B; end //??
            4'b0110:begin F=A<B; end    //A<B?F=1???F=0
            4'b0111:begin F=B<<A; end   //?B??A?
        endcase
        ZF = F==0;//F??0??ZF=1
        CF = C; //??????
        OF = A[SIZE]^B[SIZE]^F[SIZE]^C;//??????
        SF = F[SIZE];//????,?F????
        PF = ~^F;//?????F????1??F=1????1??F=0
    end     
endmodule
